module comp (input logic [7:0] a, b, output y);
    assign y = ( a == b);
endmodule
